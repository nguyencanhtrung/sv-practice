/* -------------------------------------------
* Author:   Nguyen Canh Trung
* Email:    nguyencanhtrung@me.com
* Date:     2023-09-07 08:59:19
* Filename: packages
* Last Modified by:     Nguyen Canh Trung
* Last Modified time:   2023-09-07 08:59:19
* --------------------------------------------*/
